`ifndef __UMI_OPCODES_VH__
`define __UMI_OPCODES_VH__

`define UMI_INVALID        8'b00000000
`define UMI_WRITE_NORMAL   8'b00000001
`define UMI_WRITE_RESPONSE 8'b00000010
`define UMI_WRITE_SIGNAL   8'b00000011
`define UMI_WRITE_STREAM   8'b00000100
`define UMI_WRITE_ACK      8'b00000101
`define UMI_READ           8'b00001000
`define UMI_ATOMIC_SWAP    8'b00001001
`define UMI_ATOMIC_ADD     8'b00011001
`define UMI_ATOMIC_AND     8'b00101001
`define UMI_ATOMIC_OR      8'b00111001
`define UMI_ATOMIC_XOR     8'b01001001
`define UMI_ATOMIC_MAX     8'b01011001
`define UMI_ATOMIC_MIN     8'b01101001
`define UMI_ATOMIC_USER    8'b10001001
`define UMI_USER           8'b11111111

`endif // __UMI_OPCODES_VH__
