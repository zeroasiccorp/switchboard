// Copyright (c) 2023 Zero ASIC Corporation
// This code is licensed under Apache License 2.0 (see LICENSE for details)

localparam [63:0] HEAD_OFFSET = 64'd0;
localparam [63:0] TAIL_OFFSET = 64'd64;
localparam [63:0] PACKET_OFFSET = 64'd128;
localparam PACKET_SIZE = 64;
