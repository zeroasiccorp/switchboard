* RC circuit

* Copyright (c) 2024 Zero ASIC Corporation
* This code is licensed under Apache License 2.0 (see LICENSE for details)

.SUBCKT rc in out

Rin in out 10k
Cout out 0 10p

.ENDS
