RC circuit

* Copyright (c) 2024 Zero ASIC Corporation
* This code is licensed under Apache License 2.0 (see LICENSE for details)

* voltage input
YDAC DAC0 in 0 simpleDAC
.model simpleDAC DAC (tr=5e-9 tf=5e-9)

Rin in out 10k
Cout out 0 10p

* voltage output
.measure tran ADC0 EQN V(out)

.TRAN 0 1

.END
